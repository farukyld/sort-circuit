module sort_circuit.v (
);

endmodule
